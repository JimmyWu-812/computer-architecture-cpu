module ALU_Control
(
    funct_i    (),
    ALUOp_i    (),
    ALUCtrl_o  ()
);

input [9:0] funct_i;
input [1:0] ALUOp_i;
output [2:0] ALUCtrl_o;



endmodule
